library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity controlrom is
  port (clk: in std_logic;
        addr: in std_logic_vector(8-1 downto 0);
        data: out std_logic_vector(32-1 downto 0));
end controlrom;

architecture behavioral of controlrom is
  type rom_type is array (0 to 255) of
	std_logic_vector (32-1 downto 0);

  signal ROM: rom_type := (
    "00000000000000000010000000000000",
    "00000000000010000000100000000000",
    "00000000000000010001000000000000",
    "00000000000000010001000000000001",
    "00000000000000010001000000000010",
    "00000000000000010001000000000011",
    "00000000000000010001000000000100",
    "00000000000000010001000000000101",
    "00000000000000010001000000000110",
    "00000000000000010001000000000111",
    "00000000000000010001000000001000",
    "00000000000000010001000000001001",
    "00000000000000010001000000001010",
    "00000000000000010001000000001011",
    "00000000000000010001000000001100",
    "00000000000000010001000000001101",
    "00000000000000010001000000001110",
    "00000000000000010001000000001111",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000010000010100000000110001",
    "00000000010000010100000110110000",
    "00000000010000010000000000110000",
    "00000000010000010000000000110001",
    "00000000000000000001100000000000",
    "00000000000000000100000000000000",
    "00000000000000000100000000100000",
    "00000000000000000100000000000000",
    "00000000000000000100000000000000",
    "00000000010000010000000000110001",
    "00000000000000000001000110000000",
    "00000000000000011001000000000000",
    "00000000010000010000000000100101",
    "00000000010000010000000000001010",
    "00000000000000000001000100000000",
    "00000000000100000000000101000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000001000110000000",
    "00000000000100000000000111000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000010001100000010000",
    "00000000000000010001100000010001",
    "00000000000000010001100000010010",
    "00000000000000010001100000010011",
    "00000000000000010001100000010100",
    "00000000000000010001100000010101",
    "00000000000000010001100000010110",
    "00000000000000010001100000010111",
    "00000000000000010001100000011000",
    "00000000000000010001100000011001",
    "00000000000000010001100000011011",
    "00000000000000010001100000011100",
    "00000000000000010001100000011101",
    "00000000000000010001100000011110",
    "00000000000000010001100000011111",
    "00000000000001110001000000000000",
    "00000000000001110001000000000001",
    "00000000000000000000000000000001",
    "00000000000000000000000000000001",
    "00000000000000100000000000000001",
    "00000000000000100000000000000001",
    "00000000000001000000000000000001",
    "00000000000001000000000000000001",
    "00000000000000000000000000100001",
    "00000000000000000000000000100001",
    "00000000000000100000000000100001",
    "00000000000000100000000000100001",
    "00000000000001000000000000100001",
    "00000000000001000000000000100001",
    "00000000000000000000000000000001",
    "00000000000000000000000000000001",
    "00000000000000100000000000000001",
    "00000000000000100000000000000001",
    "00000000000001000000000000000001",
    "00000000000001000000000000000001",
    "00000000000000000000000000100001",
    "00000000000000000000000000100001",
    "00000000000000100000000000100001",
    "00000000000000100000000000100001",
    "00000000000001000000000000100001",
    "00000000000001000000000000100001",
    "00000000000000000000100000000000",
    "00000000000000000000101111000000",
    "00000000000000000001100010000000",
    "00000000000100000000100011000000",
    "00000000000000000001100100010000",
    "00000000000100000000100101010000",
    "00000000000100000000000111000000",
    "00000000010000010000000000110000",
    "00000000010000010000000000110000",
    "00000000000000000000100000000000",
    "00000000000000000000101000000000",
    "00000000000000000000110000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000");

  attribute rom_style: string;
  attribute rom_style of ROM: signal is "block";

  begin
    process (addr)
    begin
        data <= ROM(conv_integer(addr));
    end process;
end behavioral;
