library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity decisionrom is
  port (clk: in std_logic;
        addr: in std_logic_vector(8-1 downto 0);
        data: out std_logic_vector(16-1 downto 0));
end decisionrom;

architecture behavioral of decisionrom is
  type rom_type is array (0 to 255) of
	std_logic_vector (16-1 downto 0);

  signal ROM: rom_type := (
    "0000000100000001",
    "0000001000000010",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "1000001010000010",
    "1000001110000011",
    "1000010010000100",
    "1000010110000101",
    "1000011010000110",
    "1000011110000111",
    "1000100010001000",
    "1000100110001001",
    "1000101010001010",
    "1000101110001011",
    "1000110010001100",
    "1000110110001101",
    "1000111010001110",
    "1000111110001111",
    "1001000010010000",
    "1001000110010001",
    "1001001010010010",
    "1001001110010011",
    "1001010010010100",
    "1001010110010101",
    "1001011010010110",
    "1001011110010111",
    "1001100010011000",
    "1001100110011001",
    "1001101010011010",
    "1001101110011011",
    "1001110010011100",
    "1001110110011101",
    "1001111010011110",
    "1011010110110101",
    "1001111110011111",
    "1010000010100000",
    "1010000110100001",
    "1010001010100010",
    "1010001110100011",
    "1010010010100100",
    "1010010110100101",
    "1010011010100110",
    "1010011110100111",
    "1010100010101000",
    "1010100110101001",
    "1010101010101010",
    "1011011010110110",
    "1010101110101011",
    "1011010110110101",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "1010110110101101",
    "1010111010101110",
    "1010111110101111",
    "1011000010110000",
    "1011000110110001",
    "1011001010110010",
    "0000000000000000",
    "0000000000000000",
    "1011001110110011",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0100111001001110",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "1011011010110100",
    "1011011010110100",
    "1011010110110100",
    "1011010010110101",
    "1011010010110101",
    "1011010110110100",
    "1011010110110100",
    "1011010010110101",
    "1011010110110100",
    "1011010010110101",
    "1011010010110101",
    "1011010110110100",
    "1011010110110100",
    "1011010010110101",
    "1011011010110100",
    "1011010010110110",
    "1011010010110110",
    "1011011010110100",
    "1011011010110100",
    "1011010010110110",
    "1011011010110100",
    "1011010010110110",
    "1011010010110110",
    "1011011010110100",
    "1011011010110100",
    "1011010010110110",
    "1010110010101100",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000");

  attribute rom_style: string;
  attribute rom_style of ROM: signal is "block";

  begin
    process (addr)
    begin
        data <= ROM(conv_integer(addr));
    end process;
end behavioral;
