library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity mainrom is
  port (clk: in std_logic;
        addr: in std_logic_vector(14-1 downto 0);
        data: out std_logic_vector(16-1 downto 0));
end mainrom;

architecture behavioral of mainrom is
  type rom_type is array (0 to 188) of
	std_logic_vector (16-1 downto 0);

  signal ROM: rom_type := (
    "0111111000000111",
    "0111111111111111",
    "0111111000000010",
    "0000000001100001",
    "0111011000111000",
    "0000000000101010",
    "0111111000000010",
    "0000110001000110",
    "0111011000111000",
    "0000000001000101",
    "0111111000000010",
    "0000000010001100",
    "0111011000111000",
    "0000000000101010",
    "0111111000000010",
    "0000000000010111",
    "0111011000111000",
    "0000000001000101",
    "0111111000000010",
    "0000000010001100",
    "0111011000111000",
    "0000000000101010",
    "0111111000000010",
    "0000000000010111",
    "0010000000010010",
    "0000110001000110",
    "0111011000111000",
    "0000000001000101",
    "0111111000000010",
    "0000000010001100",
    "0111011000111000",
    "0000000000101010",
    "0111111000000010",
    "0000000010001111",
    "0111011000111000",
    "0000000000101010",
    "0111011000111000",
    "0000000000111100",
    "0111011000111000",
    "0000000000110011",
    "0101101000000000",
    "0000000000100100",
    "1001101000010001",
    "0110100000001000",
    "0000000000000110",
    "0111011000111000",
    "0000000000110011",
    "0111101000010000",
    "0111010000000000",
    "1111111111111001",
    "0111100000111000",
    "1000000000000000",
    "1100000000000010",
    "0010101000000000",
    "0000000000000010",
    "0110100000000000",
    "1111111111111011",
    "1000001000000001",
    "1100000000000001",
    "0111100000111000",
    "1000000000000000",
    "1100000000000010",
    "0010101000000000",
    "0000000000000100",
    "0110100000000000",
    "1111111111111011",
    "1000000000000001",
    "1100000000000000",
    "0111100000111000",
    "0111111000000011",
    "0000000000000000",
    "1000100000111011",
    "0111001000010000",
    "0000000000000111",
    "0111111000000001",
    "0000000000101101",
    "0111011000111000",
    "0000000000110011",
    "0010010000010010",
    "1111111111111111",
    "0010100000010001",
    "0000000000001010",
    "0010000000001001",
    "0000000000110000",
    "1000100000111001",
    "0010011000010010",
    "0000000000001010",
    "0110110000010000",
    "1111111111111000",
    "1000101000111001",
    "0110100000001000",
    "0000000000000101",
    "0111011000111000",
    "0000000000110011",
    "0111010000000000",
    "1111111111111010",
    "0111100000111000",
    "0000000001001000",
    "0000000001100101",
    "0000000001110010",
    "0000000001100101",
    "0000000000100000",
    "0000000001100001",
    "0000000001110010",
    "0000000001100101",
    "0000000000100000",
    "0000000001110100",
    "0000000001110111",
    "0000000001101111",
    "0000000000100000",
    "0000000001101110",
    "0000000001110101",
    "0000000001101101",
    "0000000001100010",
    "0000000001100101",
    "0000000001110010",
    "0000000001110011",
    "0000000000100000",
    "0000000001100110",
    "0000000001101111",
    "0000000001101100",
    "0000000001101100",
    "0000000001101111",
    "0000000001110111",
    "0000000001100101",
    "0000000001100100",
    "0000000000100000",
    "0000000001100010",
    "0000000001111001",
    "0000000000100000",
    "0000000001110100",
    "0000000001101000",
    "0000000001100101",
    "0000000001101001",
    "0000000001110010",
    "0000000000100000",
    "0000000001110011",
    "0000000001110101",
    "0000000001101101",
    "0000000000111010",
    "0000000000001101",
    "0000000000001010",
    "0000000000000000",
    "0000000001001110",
    "0000000001101111",
    "0000000001110111",
    "0000000000100000",
    "0000000001110100",
    "0000000001111001",
    "0000000001110000",
    "0000000001100101",
    "0000000000100000",
    "0000000001110011",
    "0000000001101111",
    "0000000001101101",
    "0000000001100101",
    "0000000001110100",
    "0000000001101000",
    "0000000001101001",
    "0000000001101110",
    "0000000001100111",
    "0000000000100000",
    "0000000001100001",
    "0000000001101110",
    "0000000001100100",
    "0000000000100000",
    "0000000001001001",
    "0000000000100000",
    "0000000001110111",
    "0000000001101001",
    "0000000001101100",
    "0000000001101100",
    "0000000000100000",
    "0000000001100101",
    "0000000001100011",
    "0000000001101000",
    "0000000001101111",
    "0000000000100000",
    "0000000001101001",
    "0000000001110100",
    "0000000000100000",
    "0000000001100010",
    "0000000001100001",
    "0000000001100011",
    "0000000001101011",
    "0000000000101110",
    "0000000000001101",
    "0000000000001010",
    "0000000000000000");

  attribute rom_style: string;
  attribute rom_style of ROM: signal is "block";

  begin
    process (addr)
    begin
      if (addr <= 188) then
	data <= ROM(conv_integer(addr));
      else
	data <= (others => '0');
      end if;
    end process;
end behavioral;
